// sdram.v

// Generated using ACDS version 18.1 646

`timescale 1 ps / 1 ps
module sdram (
		input  wire        clk_clk,          //   clk.clk
		input  wire        reset_reset_n,    // reset.reset_n
		input  wire [21:0] s1_address,       //    s1.address
		input  wire [1:0]  s1_byteenable_n,  //      .byteenable_n
		input  wire        s1_chipselect,    //      .chipselect
		input  wire [15:0] s1_writedata,     //      .writedata
		input  wire        s1_read_n,        //      .read_n
		input  wire        s1_write_n,       //      .write_n
		output wire [15:0] s1_readdata,      //      .readdata
		output wire        s1_readdatavalid, //      .readdatavalid
		output wire        s1_waitrequest,   //      .waitrequest
		output wire [11:0] wire_addr,        //  wire.addr
		output wire [1:0]  wire_ba,          //      .ba
		output wire        wire_cas_n,       //      .cas_n
		output wire        wire_cke,         //      .cke
		output wire        wire_cs_n,        //      .cs_n
		inout  wire [15:0] wire_dq,          //      .dq
		output wire [1:0]  wire_dqm,         //      .dqm
		output wire        wire_ras_n,       //      .ras_n
		output wire        wire_we_n         //      .we_n
	);

	sdram_new_sdram_controller_0 new_sdram_controller_0 (
		.clk            (clk_clk),          //   clk.clk
		.reset_n        (reset_reset_n),    // reset.reset_n
		.az_addr        (s1_address),       //    s1.address
		.az_be_n        (s1_byteenable_n),  //      .byteenable_n
		.az_cs          (s1_chipselect),    //      .chipselect
		.az_data        (s1_writedata),     //      .writedata
		.az_rd_n        (s1_read_n),        //      .read_n
		.az_wr_n        (s1_write_n),       //      .write_n
		.za_data        (s1_readdata),      //      .readdata
		.za_valid       (s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (s1_waitrequest),   //      .waitrequest
		.zs_addr        (wire_addr),        //  wire.export
		.zs_ba          (wire_ba),          //      .export
		.zs_cas_n       (wire_cas_n),       //      .export
		.zs_cke         (wire_cke),         //      .export
		.zs_cs_n        (wire_cs_n),        //      .export
		.zs_dq          (wire_dq),          //      .export
		.zs_dqm         (wire_dqm),         //      .export
		.zs_ras_n       (wire_ras_n),       //      .export
		.zs_we_n        (wire_we_n)         //      .export
	);

endmodule
