`timescale 1 ps / 1 ps

module top
	(
		input 	CLK_10M,
		input		ENC_ABS_HOME,
		input 	ENC_360,
		input 	HDMI_RGB[2:0][7:0],
		output 	reg LAT,
		output 	reg SCLK,
		output 	GSCLK,
		output   SDO[11:0][3:0]

		//////////// SDRAM //////////
		output		    [12:0]		DRAM_ADDR, //address
		output		     [1:0]		DRAM_BA, //bank address
		output		          		DRAM_CAS_N, //column address strobe
		output		          		DRAM_CKE, //clock enable
		output		          		DRAM_CLK, //clock
		output		          		DRAM_CS_N, //chip select
		inout 		    [15:0]		DRAM_DQ, //SDRAM data
		output		     [1:0]		DRAM_DQM, //SDRAM byte data mask
		output		          		DRAM_RAS_N, //row address strobe
		output		          		DRAM_WE_N, //write enable
	);
	
	Pll pll(
		.clk_in_clk(CLK_10M),  			//  clk_in.clk
		.gsclk_clk(GSCLK),     			//   gsclk.clk
		.sclk_x2_clk(spiClk)    		// sclk_x2.clk // unused
	);
	
	HDMI hdmi(
		//takes the 24 HDMI_RGB values as input (they also input into top)
		//places the HDMI RGB values into SDRAM
		//we just index through SDRAM and fill it with entire 1440x720 frame
		//once it is fully populated, we switch to populating the other buffer
		//and notify the led driver code that it can start reading from memory
	);
	
	//Reading from and writing to SDRAM
	//there are 4 banks available to us
	//can we populate one bank with data while reading data from another bank
	
	
	// HDMI
	//takes in 24 bit value from HDMI decoder
	//places this information in a latch/reg to send to LED CTL
	//recieve 1440 RGB values sets for one update
	//12 by 4 by 30 by 3 array that stores the values 
	//LED CTL can assemble a length 769 bitstream from this

	// state: when finish data upload. turn off sclk
	
	//MatrixLocation
	//the spot in the matrix corresponds to the LED that the HDMI data is for

	// Reset reset(
	// 	.clk(CLK_10M),
	// 	.nReset
	// );
	
	localparam LATCH_SIZE = 'd769;
	integer bit_num = LATCH_SIZE - 1;
	reg [LATCH_SIZE:0] control_data = 769'b1100101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111000000000001010000101000010100001010000101000010100001010000101000010100001010000101000010100001010000101000010100001010000101000010100001010000101000010100001010000101000010100001010000101000010100001010000101000010100001010000101000010100001010000101000010100001010000101000010100001010000101000010100001010000101000010100001010000101000010100;
	// reg [LATCH_SIZE:0] control_data = 'b1100101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111000000000001010000101000010100001010000101000010100001010000101000010100001010000101000010100001010000101000010100001010000101000010100001010000101000010100001010000101000010100001010000101000010100001010000101000010100001010000101000010100001010000101000010100001010000101000010100001010000101000010100001010000101000010100001010000101000010100;
	
	// raw stream from arduino
	// reg [LATCH_SIZE:0] grayscale_data = 769'b0000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111;
	
	// shoving all 1's
	reg [LATCH_SIZE:0] grayscale_data = 769'b0111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
	
	// all blue
	//reg [LATCH_SIZE:0] grayscale_data = 769'b0111111111111111100000000000000000000000000000000111111111111111100000000000000000000000000000000111111111111111100000000000000000000000000000000111111111111111100000000000000000000000000000000111111111111111100000000000000000000000000000000111111111111111100000000000000000000000000000000111111111111111100000000000000000000000000000000111111111111111100000000000000000000000000000000111111111111111100000000000000000000000000000000111111111111111100000000000000000000000000000000111111111111111100000000000000000000000000000000111111111111111100000000000000000000000000000000111111111111111100000000000000000000000000000000111111111111111100000000000000000000000000000000111111111111111100000000000000000000000000000000111111111111111100000000000000000000000000000000;
	
	// all green 
	//reg [LATCH_SIZE:0] grayscale_data = 769'b0000000000000000011111111111111110000000000000000000000000000000011111111111111110000000000000000000000000000000011111111111111110000000000000000000000000000000011111111111111110000000000000000000000000000000011111111111111110000000000000000000000000000000011111111111111110000000000000000000000000000000011111111111111110000000000000000000000000000000011111111111111110000000000000000000000000000000011111111111111110000000000000000000000000000000011111111111111110000000000000000000000000000000011111111111111110000000000000000000000000000000011111111111111110000000000000000000000000000000011111111111111110000000000000000000000000000000011111111111111110000000000000000000000000000000011111111111111110000000000000000000000000000000011111111111111110000000000000000;
	
	// all red
	 //reg [LATCH_SIZE:0] grayscale_data = 769'b0000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111;

	

	reg [3:0] state = 4'd0;
	reg [30:0] iterations = 'd10;
	reg [5:0] dot_correction = 6'd127;

	
	always@(posedge CLK_10M) begin
		if (!nReset) begin
			state <= 4'd0; // initialize
			LAT <= '0;
			SCLK <= '0;
			bit_num <= LATCH_SIZE;
		end else begin
			case (state)
				4d'0: //reset all data bits to 0
					begin
						SCLK <= '0;
						data[LATCH_SIZE:0] <= '0;
					end
				4d'1: // update the data with the control data latch 
					begin
						data[768] <= '1;
						data[]
					end
			endcase

		end 
	// 	// if (!nReset) begin
	// 	// 	state <= 4'd0; // initialize
	// 	// 	LAT <= '0;
	// 	// 	SCLK <= '0;
	// 	// 	bit_num <= LATCH_SIZE;
	// 	// end else begin
	// 		case (state)
	// 			4'd9: // reset iterations
	// 				begin
	// 					iterations <= 'd10;
	// 					state <= 4'd0;
	// 				end
	// 			4'd0: // initialize, load (begin)
	// 				begin
	// 					SCLK <= '0;
	// 					if (bit_num != '0) begin							
	// 						SDO[11][3] <= (control_data >> (bit_num-1)) & 1'b1; // control_data[bit_num-1];
	// 						SDO[11][2] <= (control_data >> (bit_num-1)) & 1'b1; // control_data[bit_num-1];
	// 						SDO[11][1] <= (control_data >> (bit_num-1)) & 1'b1; // control_data[bit_num-1];
	// 						SDO[11][0] <= (control_data >> (bit_num-1)) & 1'b1; // control_data[bit_num-1];
	// 						state <= 4'd1; // initialize, shift in
	// 					end else begin
	// 						state <= 4'd2; // initialize, latch
	// 					end
	// 				end
	// 			4'd1: // initialize, shift in
	// 				begin
	// 					bit_num <= bit_num - 1;
	// 					SCLK <= '1;
	// 					state <= 4'd0; // initialize, load
	// 				end
	// 			4'd2: // initialize, latch (end)
	// 				begin
	// 					LAT <= '1;
	// 					bit_num <= LATCH_SIZE;
	// 					state <= 4'd3; // grayscale, reinit
	// 				end
	// 			4'd3: // grayscale, reinit (begin)
	// 				begin
	// 					LAT <= '0;
	// 					SCLK <= '0;
	// 					bit_num <= LATCH_SIZE;
	// 					// reset state to push control latches again after 50e6 iteratins
	// 					if (iterations == '0) begin
	// 						state <= 4'd9;
	// 					end else begin
	// 						iterations <= iterations - 1;
	// 						state <= 4'd4; // 4'd8
	// 					end
	// 				end
				
	// 			// 4'd8: // grayscale, load 0's
	// 			// 	begin
	// 			// 		SCLK <= 0;
	// 			// 		SDO[0] <= 0;
	// 			// 		SDO[1] <= 0;
	// 			// 		SDO[2] <= 0;
	// 			// 		SDO[3] <= 0;
	// 			// 		state <= 4'd5; // grayscale, shift in
	// 			// 	end
	// 			4'd4: // grayscale, load
	// 				begin
	// 					SCLK <= 0;
	// 					if (bit_num != 0) begin
	// 						SDO[11][3] <= grayscale_data[bit_num-1];
	// 						SDO[11][2] <= grayscale_data[bit_num-1];
	// 						SDO[11][1] <= grayscale_data[bit_num-1];
	// 						SDO[11][0] <= grayscale_data[bit_num-1];
	// 						state <= 4'd5; // grayscale, shift in
	// 					end else begin
	// 						state <= 4'd6; // grayscale, latch
	// 					end
	// 				end

	// 			// 4'd4: // grayscale, load 1's
	// 			// 	begin
	// 			// 		SCLK <= 0;
	// 			// 		if (bit_num != 0) begin // offset by 1 for MSB 0
	// 			// 			SDO[0] <= 1;
	// 			// 			SDO[1] <= 1;
	// 			// 			SDO[2] <= 1;
	// 			// 			SDO[3] <= 1;
	// 			// 			state <= 4'd5; // grayscale, shift
	// 			// 		end else begin
	// 			// 			state <= 4'd6; // grayscale, latch
	// 			// 		end
	// 			// 	end
				
	// 			4'd5: // grayscale, shift in
	// 				begin
	// 					bit_num = bit_num - 1;
	// 					SCLK <= '1;
	// 					state <= 4'd4; // grayscale, load
	// 				end
	// 			4'd6: // grayscale, latch (end)
	// 				begin
	// 					LAT <= '1;
	// 					bit_num <= LATCH_SIZE;
	// 					state <= 4'd3; // grayscale, reinit
	// 				end
	// 			// 4'd7: // hold loop, turn off LEDs
	// 			// 	begin
	// 			// 		LAT <= '1; // should not wipe shift register
	// 			// 		state <= 4'd7;
	// 			// 	end
	// 			default:
	// 				state <= 4'd9;
	// 		endcase
	// 	// end
	// end
endmodule